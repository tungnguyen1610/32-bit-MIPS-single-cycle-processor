package testbench_pkg;
	import uvm_pkg::*;
`include "uvm_macros.svh"
`include "sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "agent.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "subscriber.sv"
`include "env.sv"
`include "test.sv"


endpackage : testbench_pkg   // <-- must be present
